module states(input CLK,
	      input 	       RST,
	      input 	       CHANGE_REQUESTED,
	      input [2:0]      COMMAND,
	      output 	       CHANGE_POSSIBLE,
	      output reg [2:0] STATE,
	      output reg       CLOCK_COMMAND);
  reg [1:0] 	     counter;
  reg 		     state_is_readwrite;

  assign CHANGE_POSSIBLE = ((counter == 2'h3) ||
			    (state_is_readwrite && (COMMAND == STATE))) ?
			   1 : 0;

  always @(posedge CLK)
    if (!RST)
      begin
	counter <= 2'h3;
	state_is_readwrite <= 0;
	CLOCK_COMMAND <= 1'b0;
	STATE <= `PRCH;
      end
    else
      if (CHANGE_POSSIBLE)
	begin
	  if (CHANGE_REQUESTED)
	    begin
	      STATE <= COMMAND;
	      state_is_readwrite <= ((COMMAND == `READ) || (COMMAND == `WRTE));

	      if (COMMAND == `ACTV)
		counter <= 2'h1;
	      else
		counter <= 2'h0;

	      if (COMMAND == `PRCH)
		CLOCK_COMMAND <= 1'b1;
	      else
		CLOCK_COMMAND <= 1'b0;
	    end
	end // if (CHANGE_POSSIBLE)
      else
	begin
	  CLOCK_COMMAND <= 1'b0;

	  if ((CHANGE_REQUESTED & state_is_readwrite) && (COMMAND == STATE))
	    counter <= 2'h0;
	  else
	    counter <= counter +1;
	end

endmodule // states

module enter_state(input CLK,
		   input 	    RST,
		   input [11:0]     PAGE_REQUEST,
		   input 	    WE,
		   input 	    DO_ACT,
		   input 	    CHANGE_POSSIBLE,
		   input 	    CLOCK_COMMAND,
		   output reg [2:0] COMMAND,
		   output 	    CHANGE_REQUESTED,
		   output 	    DO_WRITE);
  reg [11:0] 			    page_current;
  reg [2:0] 			    command_sequence[2:0];
  reg [1:0] 			    command_len;
  reg 				    we_sequence[2:0];

  wire [2:0] 			    rw_command;

  assign CHANGE_REQUESTED = (command_len == 2'h3) ? 0 : 1;
  assign rw_command = WE ? `WRTE : `READ;
  assign DO_WRITE = we_sequence[command_len];

  always @(posedge CLK)
    if (!RST)
      begin
	page_current <= 0; /* TODO: will have to be hacked */
	command_sequence <= {`NOP/*actually PRCH*/,`ACTV,`READ};
	command_len <= 2'h3;
	COMMAND <= `NOP;
      end
    else
      begin
	if (CHANGE_REQUESTED)
	  begin
	    if (CHANGE_POSSIBLE)
	      begin
		command_len <= command_len +1;
		COMMAND <= command_sequence[command_len];
		page_current <= PAGE_REQUEST;
		/* TODO: setup data receivers/senders here */
	      end
	    else
	      if (CLOCK_COMMAND)
		COMMAND <= `PRCH;
	      else
		COMMAND <= `NOP;
	  end // if (CHANGE_REQUESTED)
	else
	  begin
	    command_sequence <= {`NOP/*actually PRCH*/,`ACTV,rw_command};
	    we_sequence <= {1'b0,1'b0,WE};

	    if (DO_ACT)
	      begin
		if (PAGE_REQUEST == page_current)
		  command_len <= 2'h2;
		else
		  command_len <= 2'h0;
	      end
	  end // else: !if(CHANGE_REQUESTED)
      end

endmodule // enter_state

module outputs(input CLK_p,
	       input 		 CLK_n,
	       input 		 CLK_d,
	       input 		 RST,
	       input 		 CHANGE_REQUESTED,
	       input 		 CHANGE_POSSIBLE,
	       input [31:0] 	 DATA_W,
	       input 		 WE,
	       inout [15:0] 	 DQ,
	       inout 		 DQS,
	       output reg [31:0] DATA_R,
	       output reg 	 DATA_VALID);
  reg [15:0] 			 dq_driver;
  reg [31:0] 			 dq_driver_pre, dq_driver_holdlong;
  reg 				 dqs_driver, pipe_clk_dqs;
  reg 				 will_write, do_write, do_deltawrite, do_halfwrite;
  reg 				 will_read, really_will_read, about_to_read,
				 do_read, reading;

  assign DQ = do_deltawrite ? dq_driver : {{16}1'bz};
  assign DQS = (do_write | do_halfwrite) ? dqs_driver : 1'bz;

  always @(CLK_n)
    dqs_driver <= CLK_n;

  always @(posedge CLK_n)
    if (!RST)
      begin
	dq_driver_pre <= 0;
	will_read <= 0;
	will_write <= 0;
	do_read <= 0;
	about_to_read <= 0;
	really_will_read <= 0;
	do_write <= 0;
	dq_driver_holdlong <= 0;
      end
    else
      begin
	will_write <= 0;
	do_write <= will_write;
	dq_driver_holdlong <= dq_driver_pre;

	will_read <= 0;
	really_will_read <= will_read;
	about_to_read <= really_will_read;
	do_read <= about_to_read;

	if (CHANGE_REQUESTED & CHANGE_POSSIBLE)
	  begin
	    if (WE)
	      begin
		will_write <= 1;
	      end
	    else
	      will_read <= 1;

	    dq_driver_pre <= DATA_W;
	  end // if (CHANGE_REQUESTED & CHANGE_POSSIBLE)
      end // else: !if(!RST)

  always @(posedge CLK_p)
    if (!RST)
      begin
	do_halfwrite <= 0;
	reading <= 0;
      end
    else
      begin
	do_halfwrite <= do_write;
	reading <= do_read;
      end

  always @(CLK_d)
    if (!RST)
      begin
	do_deltawrite <= 0;
	dq_driver <= 0;
	DATA_R <= 0;
	DATA_VALID <= 0;
      end
    else
      begin
	do_deltawrite <= do_write;

	if (dqs_driver)
	  begin
	    dq_driver <= dq_driver_holdlong[15:0];
	    DATA_R[31:16] <= DQ;
	  end
	else
	  begin
	    dq_driver <= dq_driver_holdlong[31:16];
	    DATA_R[15:0] <= DQ;
	    DATA_VALID <= reading;
	  end
      end

endmodule // outputs
